 module Tb0000000001 ();
 reg clk_in;
 reg clk_out;
 reg rst;
 wire data_in;
 reg data_valid;
 wire data_out;
 reg [31:0] tx_data_buffer;
 reg data_in_reg;
 wire is_frame_sychronized;
 wire [2:0] synchronizer_state;
 wire data_sync_out;
 wire data_decoder_out;
 initial begin
    clk_in = 0;
    clk_out = 1;
 end
 always #10 clk_in = ~clk_in;  // 20ns����
 always #5 clk_out = ~clk_out; // 10ns����
 assign data_in = data_in_reg;
 // Instantiate the Hamming Encoder
HammingEncoder0000000001  u_0000000001_HammingEncoder0000000001(.clk_in(clk_in), .clk_out(clk_out), .rst(rst), .data_in(data_in), .data_valid(data_valid), .data_out(data_out), .data_in_ready(data_in_ready));
 // Instantiate frame synchronizer
SyncFrame0000000001  u_0000000001_SyncFrame0000000001(.clk_out(clk_out), .rst(rst), .data_in(data_out), .is_frame_sychronized(is_frame_sychronized), .synchronizer_state(synchronizer_state), .data_sync_out(data_sync_out));
 // Instantiate the Hamming Decoder
Decoder0000000001  u_0000000001_Decoder0000000001(.clk_decoder_in(clk_out), .clk_decoder_out(clk_in), .rst(rst), .decoder_data_valid(is_frame_sychronized), .data_decoder_in(data_sync_out), .data_decoder_out(data_decoder_out));
 task send_data;
     input [31:0] data;
     integer i;
     begin
         for (i = 31; i >= 0; i = i - 1) begin
             data_in_reg = data[i];
             data_valid = 1;
             @(posedge clk_in);
         end
         data_valid = 0;
     end
 endtask
 initial begin
     $dumpfile("wave.vcd");
     $dumpvars(0, Tb0000000001);
     # 5
     rst = 1'b1;
     # 20 rst = 1'b0;
     # 20 data_valid = 1'b1;
     @ (posedge clk_in);
     send_data(32'b00000000011111001100110101111101);
     send_data(32'b10001101010111100111101101101010);
     send_data(32'b01010011011111100011000110011111);
     send_data(32'b01001110010001001001011100101101);
     send_data(32'b11111001100001101101011110001111);
     send_data(32'b01110000110100110001010111101010);
     send_data(32'b11101101011011011011101001010101);
     send_data(32'b10001111001101100010111110100100);
     send_data(32'b00111110111010000110110110010011);
     send_data(32'b01000000111100111111101010110001);
     send_data(32'b10111001001000001010000100000001);
     send_data(32'b01011101001000010001110000100110);
     send_data(32'b01000110011011010000010101111101);
     send_data(32'b11001000110000001110010010111011);
     send_data(32'b11101101011010011101010101110000);
     send_data(32'b11001011110010000101111100101001);
     send_data(32'b10100011111011011110111011000111);
     send_data(32'b00101100110000011100001010001110);
     send_data(32'b10110011000111011010011000101111);
     send_data(32'b01111110100010100000100111110011);
     send_data(32'b00000111100100100100000111001010);
     send_data(32'b01110110010010111110001010110011);
     send_data(32'b10010001100111001110111000000100);
     send_data(32'b01010110000000001100110011010010);
     send_data(32'b10000010000010001111100010110000);
     send_data(32'b10100001011111100001101001101001);
     send_data(32'b11010101101001011110100011100110);
     send_data(32'b10010101011001011111111111110010);
     send_data(32'b11101100001011110000000111110001);
     send_data(32'b00110010110011110110100000000100);
     send_data(32'b10111011100010000100000110101000);
     send_data(32'b11011101011110101111100010101000);
     send_data(32'b00111001010100000011111100000000);
     send_data(32'b11110011000001101100001011010001);
     send_data(32'b10111000100010111110101110011000);
     send_data(32'b01101010110110011100110110111001);
     send_data(32'b01111010011001011111110011100101);
     send_data(32'b10110100010101000110000010011011);
     send_data(32'b10011111101010110111101001011101);
     send_data(32'b11000100010110000001100110101111);
     send_data(32'b01110001101111011001001010101011);
     send_data(32'b00010101001110011011000100100000);
     send_data(32'b11010101101100101111010001100101);
     send_data(32'b00011010101100101111010001010100);
     send_data(32'b00001100000011010010101110111100);
     send_data(32'b11111011101010011010110111110111);
     send_data(32'b01000100001010010111011110001100);
     send_data(32'b01010011011000111101101010000001);
     send_data(32'b00110011001111111100001100010111);
     send_data(32'b01000000000011000110001010001110);
     send_data(32'b00100010101110110000010101001101);
     send_data(32'b10101110101000011100110011000100);
     send_data(32'b11110010101110111000101001001110);
     send_data(32'b01111101111110100101000110000101);
     send_data(32'b00010110001100011011000010110000);
     send_data(32'b11010010010000111010010111011100);
     send_data(32'b01101011000101000100011110110001);
     send_data(32'b10110111001001001001101110011101);
     send_data(32'b11011110010110011100010101010101);
     send_data(32'b01011111100001011111010001000110);
     send_data(32'b11000111011001111011110000100111);
     send_data(32'b10111001111011111101110101010101);
     send_data(32'b00001001101110000001101001011011);
     send_data(32'b00110011111111100010111001110100);
     send_data(32'b00001011111000101011100000011010);
     send_data(32'b01111100000010101010100111010011);
     send_data(32'b10111000111101101001101100000110);
     send_data(32'b01101000000010010111101110000001);
     send_data(32'b01010001111111001100101111101001);
     send_data(32'b10011000000000101010000100000110);
     send_data(32'b00100000110010001100011111000011);
     send_data(32'b10110011111001000000101110001110);
     send_data(32'b11000101010111001100100000111110);
     send_data(32'b11001001101111010001101001010010);
     send_data(32'b00001001011010010110111000000000);
     send_data(32'b00111110111101111001111000001010);
     send_data(32'b01101110011100001001001000000111);
     send_data(32'b10110111110011101110100100010110);
     send_data(32'b01010000001011011011000010100011);
     send_data(32'b01100110001000111011001111111010);
     send_data(32'b00100010101001010101001100010001);
     send_data(32'b11100000001100011001110001111101);
     send_data(32'b11101100011011011111010011101000);
     send_data(32'b10101001010000010100110110011001);
     send_data(32'b11000000111010100011011110001111);
     send_data(32'b10000111001100000110110101010111);
     send_data(32'b00101001100111001110000100000111);
     send_data(32'b10000111110011111011000101011011);
     send_data(32'b10110101110100000010010101110111);
     send_data(32'b10001100000101101001110100011010);
     send_data(32'b01111110000001010011010011111010);
     send_data(32'b00011110011101001111000110110100);
     send_data(32'b01110011101001000000001011010111);
     send_data(32'b11000101001101001010001000100101);
     send_data(32'b01011100111001111011101101000110);
     send_data(32'b11101000101001111010101111001100);
     send_data(32'b01111111110001001010100010000010);
     send_data(32'b00010100110000011100111111000010);
     send_data(32'b11111111000101010000000110001100);
     send_data(32'b00101101111110010010000000111001);
     # 1500 $finish;
 end
 integer fd;
 integer fd_decoder_out;
 initial begin
   fd = $fopen("encoded_bits.txt", "w");
   fd_decoder_out = $fopen("decoder_out_bits.txt", "w");
 end
 always @(posedge clk_out) begin
   // $display("Time:%t Output bit: %b", $time, data_out);
   $fdisplay(fd, "%b", data_out);
 end
 always @(posedge clk_in) begin
   $fdisplay(fd_decoder_out, "%b", data_decoder_out);
 end
 endmodule
